module top_module (
    input in,
    output out);
assign out = 1'b0;
   
endmodule