module top_module (
    input clk,
    input d, 
    input ar,   // asynchronous reset
    output q);
 wire out1,out2;
    always @(posedge clk or posedge ar) 
        begin
        if(ar==1) 
            begin
            q<=0;
        end
        else if(ar==0) begin
            q<=d;
        end
    end
endmodule
