module top_module( output zero );

// Insert your code here
    assign zero = 1'b0;

endmodule
