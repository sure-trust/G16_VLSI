module top_module (
    input d, 
    input ena,
    output q);
wire in,out1,out2;
    always @(*) begin
        out1=~(out2|(~d)&ena);
        out2=~(out1 | d&ena);
        q=out1;
    end
endmodule
