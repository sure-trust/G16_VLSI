module top_module (
    input clk,
    input x,
    output reg z
); 
	reg out1=0, out2, out3;
    initial z = 1;
    always @(posedge clk) begin
        out1 <= x ^ out1;
        out2 <= x & ~out2;
        out3 <= x | ~out3;
        z <= ~(out1 | out2 | out3);
    end
endmodule
