module top_module (
    input [3:0]clk,
    input [1:0]reset,
    input [1:0]enable,
    output [3:0] Q,
    output c_enable,//enables the clock when the reset pin goes to high state
    output c_load,//c load takes 1 bit to load the c_d
    output [3:0] c_d
  ); //
  wire [3:0] Q_tmp;
  assign c_enable=enable;
  assign c_d=c_load?1:0;
  always @(posedge clk)
  begin
    if(reset)
    begin
      Q <= 1;
      Q_tmp <= 1;
    end
    else
    begin
      if(enable)
      begin
        if(Q == 12)
        begin
          Q <= 1;
          Q_tmp <= 1;
        end
        else
        begin
          Q <= Q + 1;
          Q_tmp <= Q_tmp + 1;
        end
      end
    end
  end

  always @(*)
  begin
    if(reset || (Q == 12 && c_enable))
    begin
      c_load <= 1;
    end
    else
    begin
      c_load <= 0;
    end
  end

  count4 the_counter (clk, c_enable, c_load, c_d, Q_tmp);

endmodule
