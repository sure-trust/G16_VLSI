module top_module(input a,input b,output out);
    mod_a ins(a,b,out);
endmodule