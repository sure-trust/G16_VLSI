module top_module( 
    input a, 
    input b, 
    output out );
    nor (out,b,a);
endmodule