module top_module (
    input clk,
    input in, 
    output out);
    wire out1,out2;
    always @(posedge clk) begin
        out1=out2^in;
        out2=out1;
        out=out2;
    end
endmodule